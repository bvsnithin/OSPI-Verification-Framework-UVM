package agent_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "ospi_sequencer.sv"
  `include "ospi_driver.sv"
  `include "ospi_monitor.sv"
  `include "ospi_agent.sv"

endpackage
