

module ospi_ctrl (
    input logic        clk,
    input  logic       rst_n,
    // Interface signals connecting to the pins
    input  logic       cs_n,
    input  logic       sclk,
    inout  wire [7:0]  dq,
    inout  wire        dqs
);
    logic [7:0] mem [0:255];
    logic [7:0] data_out;
    logic       drive_bus;

    // Tri-state buffer for the Bidirectional DQ bus
    assign dq = drive_bus ? data_out : 8'bz;

    // Basic Reset Logic
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            drive_bus <= 0;
            data_out  <= 0;
        end 
        else begin
        // This is where the actual Controller logic goes.
        // For now, we leave it passive to ensure the testbench compiles.
        end
    end


endmodule: ospi_ctrl