package env_pkg;

  import uvm_pkg::*;
  import agent_pkg::*;
  `include "uvm_macros.svh"

  // `include "virtual_sequencer.sv"
  `include "ospi_scoreboard.sv"
  `include "ospi_env.sv"
  

endpackage
